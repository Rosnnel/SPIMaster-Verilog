// SPDX-License-Identifier: CERN-OHL-S-2.0
// © 2025 Rosnnel Moncada

module PISOZReg #(parameter WordLen=8)
(clk,ShiftEdge,EnPISO,LoadPISO,WordFlg,TristateMode,BitOrder,DataIN,MOSI,HBReceviedData);

    input TristateMode;
    input clk,ShiftEdge,EnPISO,LoadPISO,WordFlg,BitOrder;
    input [WordLen-1:0] DataIN;
    output [WordLen-1:0]HBReceviedData;
    inout MOSI;

    reg [WordLen-1:0] TXReg,RXReg;

    always@(posedge clk)
    begin
        if(EnPISO)
        begin
            if(TristateMode) //Transmitting Data
            begin
                if(LoadPISO)
                    TXReg <= DataIN;
                else if(ShiftEdge && ~WordFlg)
                begin
                    if(BitOrder)      //Little Endian
                        TXReg <= {1'b0,TXReg[WordLen-1:1]};
                    else                //Big Endian
                        TXReg <= {TXReg[WordLen-2:0],1'b0};
                end
            end
            else if(~TristateMode) //Receiving Data
            begin
                if(ShiftEdge && ~WordFlg)
                begin
                    if(~BitOrder)      //Little Endian
                        RXReg <= {MOSI,RXReg[WordLen-1:1]};
                    else                //Big Endian
                        RXReg <= {RXReg[WordLen-2:0],MOSI};
                end
            end
        end
    end

    assign MOSI = (TristateMode) ? ((BitOrder) ? TXReg[0] : TXReg[WordLen-1]) : 1'bz;
    assign HBReceviedData = RXReg;

endmodule